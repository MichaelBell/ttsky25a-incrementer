MACRO logo
  CLASS BLOCK ;
  FOREIGN logo ;
  ORIGIN -8.700 -7.200 ;
  SIZE 108.600 BY 106.200 ;
  OBS
      LAYER met4 ;
        RECT 8.700 7.200 117.300 113.400 ;
  END
END logo
END LIBRARY

