magic
tech sky130A
timestamp 1752183585
<< nwell >>
rect -30 -20 390 135
<< pwell >>
rect -20 -151 380 -44
<< nmos >>
rect 25 -125 40 -63
rect 125 -125 140 -63
rect 173 -125 188 -63
rect 273 -125 288 -63
rect 325 -125 340 -63
<< pmos >>
rect 25 0 40 95
rect 125 0 140 95
rect 225 0 240 95
rect 325 0 340 95
<< ndiff >>
rect -4 -125 69 -63
rect 96 -125 169 -63
rect 144 -125 217 -63
rect 244 -125 317 -63
rect 296 -125 369 -63
<< pdiff >>
rect -4 0 69 95
rect 96 0 169 95
rect 196 0 269 95
rect 296 0 369 95
<< ndiffc >>
rect 0 -115 17 -75
rect 48 -110 65 -70
rect 100 -110 117 -80
rect 148 -110 165 -90
rect 196 -115 213 -80
rect 248 -110 265 -80
rect 298 -120 317 -103
rect 348 -110 365 -80
<< pdiffc >>
rect 0 20 17 80
rect 48 20 65 80
rect 100 50 117 80
rect 148 50 165 80
rect 200 20 217 80
rect 248 20 265 80
rect 300 50 317 80
rect 348 50 365 80
<< poly >>
rect 25 -139 40 108
rect 75 -46 125 -19
rect 40 -51 125 -14
rect 125 -139 140 108
rect 173 -139 188 -14
rect 188 -51 273 -14
rect 273 -139 288 -14
rect 225 -15 240 109
rect 325 -139 340 108
rect 325 -46 362 -19
<< polycont >>
rect 85 -41 115 -24
rect 185 -41 215 -24
rect 335 -41 352 -24
<< locali >>
rect 82 -49 118 -16
rect 0 -125 17 -65
rect 0 10 17 90
rect 48 -120 65 90
rect 100 -120 117 -70
rect 148 -120 165 -80
rect 100 40 117 90
rect 148 40 165 90
rect 65 1 175 18
rect 158 -49 175 1
rect 175 -49 225 -16
rect 196 -125 213 -70
rect 248 -120 265 -70
rect 200 10 217 130
rect 248 -15 265 90
rect 325 -44 362 -21
rect 265 -15 342 2
rect 325 -21 342 -15
rect 298 -128 317 -98
rect 298 40 317 90
rect 225 -49 308 -32
rect 348 -120 365 -61
rect 291 -61 308 -49
rect 291 -78 356 -61
rect 348 40 365 90
<< viali >>
rect 0 -115 17 -75
rect 0 20 17 80
rect 82 -41 99 -24
rect 100 -110 117 -80
rect 148 -120 165 -100
rect 100 40 117 70
rect 148 50 165 80
rect 196 -115 213 -80
rect 248 -110 265 -80
rect 200 20 217 60
rect 248 20 265 60
rect 298 -120 317 -95
rect 298 50 317 80
rect 348 50 365 80
<< metal1 >>
rect -20 -167 50 -127
rect -3 -127 50 -121
rect -20 97 20 137
rect -3 86 20 97
rect -3 -121 50 -69
rect -3 14 20 86
rect 65 -47 102 -18
rect 97 -120 120 -62
rect 145 -126 168 -94
rect 97 0 120 80
rect 145 44 168 86
rect 116 -80 133 32
rect 147 -120 168 0
rect 193 -121 219 -74
rect 245 -120 271 70
rect 197 0 220 70
rect 168 -20 220 0
rect 295 -126 320 85
rect 145 85 320 105
rect 342 -53 368 86
rect 65 -140 82 -40
rect 65 -155 168 -140
<< via1 >>
rect 71 -47 97 -21
rect 342 -47 368 -21
rect 97 6 123 32
rect 245 6 271 32
rect 20 -115 46 -85
rect 193 -115 219 -85
<< metal2 >>
rect 65 -47 371 -21
rect 97 0 271 38
rect 20 -125 219 -75
<< labels >>
<< end >>
