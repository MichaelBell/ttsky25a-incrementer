MACRO logo
  CLASS BLOCK ;
  FOREIGN logo ;
  ORIGIN -8.800 -7.200 ;
  SIZE 108.400 BY 106.000 ;
  OBS
      LAYER met4 ;
        RECT 8.800 7.200 117.200 113.200 ;
  END
END logo
END LIBRARY

