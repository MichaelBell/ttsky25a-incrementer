magic
tech sky130A
timestamp 1757258261
<< metal4 >>
rect 6150 11310 6240 11340
rect 6120 11250 6270 11310
rect 6120 11220 6300 11250
rect 7170 11220 7260 11250
rect 6090 11100 6300 11220
rect 7140 11190 7290 11220
rect 7140 11160 7320 11190
rect 7110 11130 7320 11160
rect 6090 10980 6330 11100
rect 7110 11070 7350 11130
rect 7110 11040 7380 11070
rect 7080 11010 7380 11040
rect 6090 10890 6360 10980
rect 7080 10920 7410 11010
rect 6120 10800 6390 10890
rect 7080 10860 7440 10920
rect 7050 10830 7440 10860
rect 6120 10710 6420 10800
rect 6150 10680 6450 10710
rect 7050 10680 7230 10830
rect 7290 10770 7470 10830
rect 7290 10740 7500 10770
rect 7320 10710 7500 10740
rect 7320 10680 7530 10710
rect 6150 10620 6480 10680
rect 7050 10620 7200 10680
rect 7350 10650 7560 10680
rect 6150 10560 6510 10620
rect 6180 10530 6540 10560
rect 6180 10500 6570 10530
rect 6180 10410 6360 10500
rect 6390 10470 6570 10500
rect 7020 10470 7200 10620
rect 7380 10620 7560 10650
rect 7380 10590 7590 10620
rect 7410 10560 7620 10590
rect 7440 10500 7650 10560
rect 7470 10470 7680 10500
rect 6390 10440 6600 10470
rect 7020 10440 7170 10470
rect 7500 10440 7710 10470
rect 6210 10380 6360 10410
rect 6420 10380 6630 10440
rect 6210 10230 6390 10380
rect 6450 10350 6660 10380
rect 6480 10290 6690 10350
rect 6990 10320 7170 10440
rect 7530 10410 7740 10440
rect 7560 10350 7770 10410
rect 7470 10320 7800 10350
rect 6510 10260 6720 10290
rect 6240 10200 6390 10230
rect 6540 10230 6750 10260
rect 6540 10200 6780 10230
rect 6960 10200 7140 10320
rect 7440 10290 7830 10320
rect 7380 10260 7860 10290
rect 7320 10230 7620 10260
rect 7650 10230 7890 10260
rect 7260 10200 7590 10230
rect 7680 10200 7920 10230
rect 6240 9840 6420 10200
rect 6570 10170 6810 10200
rect 6600 10140 6810 10170
rect 6930 10140 7110 10200
rect 7200 10170 7560 10200
rect 7710 10170 7950 10200
rect 7170 10140 7530 10170
rect 7740 10140 7980 10170
rect 6630 10110 6840 10140
rect 6900 10110 7110 10140
rect 7140 10110 7470 10140
rect 7770 10110 8010 10140
rect 6660 10080 6870 10110
rect 6900 10080 7080 10110
rect 6660 10050 7080 10080
rect 7140 10080 7410 10110
rect 7800 10080 8040 10110
rect 7140 10050 7350 10080
rect 7830 10050 8070 10080
rect 6690 10020 7050 10050
rect 7140 10020 7290 10050
rect 7860 10020 8070 10050
rect 6720 9990 7050 10020
rect 7170 9990 7260 10020
rect 7890 9990 8100 10020
rect 6750 9960 7050 9990
rect 7890 9960 8130 9990
rect 6780 9930 7020 9960
rect 7920 9930 8160 9960
rect 6810 9900 7020 9930
rect 7950 9900 8190 9930
rect 6600 9870 6750 9900
rect 6810 9870 7050 9900
rect 7980 9870 8220 9900
rect 6570 9840 6780 9870
rect 6840 9840 7080 9870
rect 8010 9840 8250 9870
rect 6240 9780 6390 9840
rect 6510 9810 6780 9840
rect 6870 9810 7110 9840
rect 8040 9810 8250 9840
rect 6480 9780 6780 9810
rect 6900 9780 7140 9810
rect 8040 9780 8280 9810
rect 6210 9570 6390 9780
rect 6450 9750 6780 9780
rect 6930 9750 7170 9780
rect 8010 9750 8310 9780
rect 6450 9720 6750 9750
rect 6960 9720 7200 9750
rect 7980 9720 8310 9750
rect 6480 9690 6630 9720
rect 6990 9690 7230 9720
rect 7950 9690 8340 9720
rect 7020 9660 7260 9690
rect 7890 9660 8340 9690
rect 7050 9630 7290 9660
rect 7860 9630 8130 9660
rect 8160 9630 8370 9660
rect 7080 9600 7350 9630
rect 7800 9600 8100 9630
rect 7110 9570 7380 9600
rect 7590 9570 8070 9600
rect 8190 9570 8370 9630
rect 6210 9480 6360 9570
rect 7140 9540 7410 9570
rect 7560 9540 8040 9570
rect 7200 9510 7440 9540
rect 7530 9510 7980 9540
rect 7230 9480 7470 9510
rect 6180 9000 6360 9480
rect 7260 9450 7470 9480
rect 7530 9480 7920 9510
rect 7530 9450 7860 9480
rect 6930 9420 7050 9450
rect 7290 9420 7500 9450
rect 7560 9420 7770 9450
rect 6900 9390 7080 9420
rect 7320 9390 7530 9420
rect 8220 9390 8400 9570
rect 6840 9360 7080 9390
rect 7350 9360 7560 9390
rect 6600 9330 7080 9360
rect 6570 9300 7050 9330
rect 7380 9300 7590 9360
rect 6570 9270 7020 9300
rect 7410 9270 7620 9300
rect 6570 9240 6960 9270
rect 7440 9240 7650 9270
rect 6570 9210 6900 9240
rect 7470 9210 7650 9240
rect 6630 9180 6780 9210
rect 7470 9180 7680 9210
rect 7500 9150 7680 9180
rect 8250 9150 8400 9390
rect 7530 9060 7710 9150
rect 6210 8880 6360 9000
rect 7560 8970 7740 9060
rect 8220 9000 8400 9150
rect 8160 8970 8400 9000
rect 7380 8940 7500 8970
rect 7350 8910 7500 8940
rect 7290 8880 7530 8910
rect 6210 8760 6390 8880
rect 7260 8850 7530 8880
rect 7590 8850 7770 8970
rect 8130 8940 8400 8970
rect 8100 8910 8400 8940
rect 8070 8880 8370 8910
rect 8040 8850 8370 8880
rect 7200 8820 7500 8850
rect 7620 8820 7770 8850
rect 8010 8820 8370 8850
rect 6600 8790 6750 8820
rect 7110 8790 7470 8820
rect 6240 8730 6390 8760
rect 6570 8760 7410 8790
rect 6570 8730 7380 8760
rect 5640 8700 5670 8730
rect 5580 8670 5730 8700
rect 5580 8640 5760 8670
rect 5550 8610 5790 8640
rect 6240 8610 6420 8730
rect 6570 8700 7320 8730
rect 6600 8670 7260 8700
rect 6690 8640 7200 8670
rect 7620 8640 7800 8820
rect 7860 8790 8370 8820
rect 7830 8760 8370 8790
rect 7830 8730 8160 8760
rect 7830 8700 8130 8730
rect 7860 8670 8040 8700
rect 6780 8610 7080 8640
rect 7650 8610 7800 8640
rect 5550 8580 5850 8610
rect 5550 8550 5880 8580
rect 5550 8520 5940 8550
rect 6270 8520 6450 8610
rect 5520 8490 6000 8520
rect 5520 8460 5700 8490
rect 5730 8460 6060 8490
rect 6300 8460 6480 8520
rect 5520 8430 5670 8460
rect 5760 8430 6120 8460
rect 5490 8370 5670 8430
rect 5820 8400 6180 8430
rect 6330 8400 6510 8460
rect 5880 8370 6270 8400
rect 6360 8370 6540 8400
rect 5460 8280 5640 8370
rect 5940 8340 6330 8370
rect 6360 8340 6570 8370
rect 7650 8340 7830 8610
rect 5970 8310 6570 8340
rect 7680 8310 7830 8340
rect 8190 8520 8370 8760
rect 8190 8400 8340 8520
rect 6030 8280 6600 8310
rect 5430 8220 5610 8280
rect 6090 8250 6630 8280
rect 6180 8220 6630 8250
rect 7020 8220 7080 8250
rect 5400 8160 5580 8220
rect 6240 8190 6660 8220
rect 6720 8190 7320 8220
rect 6300 8160 7410 8190
rect 7680 8160 7860 8310
rect 5370 8100 5550 8160
rect 6360 8130 7500 8160
rect 6360 8100 7560 8130
rect 5340 8070 5550 8100
rect 6270 8070 7620 8100
rect 5340 8010 5520 8070
rect 6180 8040 6840 8070
rect 7170 8040 7680 8070
rect 7710 8040 7890 8160
rect 6090 8010 6660 8040
rect 7320 8010 7860 8040
rect 5310 7950 5490 8010
rect 6030 7980 6540 8010
rect 7410 7980 7800 8010
rect 5970 7950 6450 7980
rect 7500 7950 7830 7980
rect 5280 7860 5460 7950
rect 5910 7920 6360 7950
rect 7560 7920 7890 7950
rect 5850 7890 6270 7920
rect 7620 7890 7920 7920
rect 8190 7890 8370 8400
rect 5790 7860 6180 7890
rect 7650 7860 7950 7890
rect 5280 7830 5430 7860
rect 5730 7830 6120 7860
rect 7710 7830 8010 7860
rect 5250 7770 5430 7830
rect 5670 7800 6060 7830
rect 7770 7800 8040 7830
rect 5610 7770 5970 7800
rect 7800 7770 8070 7800
rect 8220 7770 8370 7890
rect 5250 7680 5400 7770
rect 5550 7740 5910 7770
rect 7830 7740 8100 7770
rect 5490 7710 5880 7740
rect 7890 7710 8130 7740
rect 5460 7680 5820 7710
rect 7920 7680 8160 7710
rect 8220 7680 8400 7770
rect 5250 7650 5760 7680
rect 7950 7650 8190 7680
rect 8250 7650 8370 7680
rect 5250 7620 5700 7650
rect 7980 7620 8220 7650
rect 8280 7620 8340 7650
rect 5250 7590 5640 7620
rect 8010 7590 8250 7620
rect 5250 7560 5580 7590
rect 8040 7560 8280 7590
rect 5250 7530 5520 7560
rect 8070 7530 8310 7560
rect 5250 7500 5490 7530
rect 8100 7500 8340 7530
rect 5250 7470 5430 7500
rect 8130 7470 8340 7500
rect 5250 7440 5370 7470
rect 8160 7440 8370 7470
rect 5250 7410 5340 7440
rect 6330 7410 6570 7440
rect 6270 7380 6660 7410
rect 8190 7380 8400 7440
rect 6240 7350 6720 7380
rect 8220 7350 8430 7380
rect 6210 7320 6780 7350
rect 8250 7320 8460 7350
rect 6180 7290 6780 7320
rect 6150 7260 6780 7290
rect 8280 7290 8460 7320
rect 8280 7260 8490 7290
rect 6120 7230 6360 7260
rect 6600 7230 6750 7260
rect 8310 7230 8490 7260
rect 6090 7200 6330 7230
rect 6660 7200 6720 7230
rect 8310 7200 8520 7230
rect 6060 7170 6300 7200
rect 8340 7170 8520 7200
rect 6060 7140 6270 7170
rect 8340 7140 8550 7170
rect 6030 7110 6240 7140
rect 6030 7080 6210 7110
rect 8370 7080 8550 7140
rect 6000 7050 6210 7080
rect 7500 7050 7530 7080
rect 6000 7020 6180 7050
rect 5970 6930 6150 7020
rect 7440 6990 7590 7050
rect 8400 7020 8580 7080
rect 7440 6930 7620 6990
rect 8430 6930 8610 7020
rect 5940 6840 6120 6930
rect 7470 6870 7650 6930
rect 8460 6870 8640 6930
rect 7500 6840 7650 6870
rect 8490 6840 8640 6870
rect 5910 6690 6090 6840
rect 7500 6780 7680 6840
rect 8490 6780 8670 6840
rect 7530 6720 7680 6780
rect 5910 6450 6060 6690
rect 5910 6210 6090 6450
rect 7530 6420 7710 6720
rect 8520 6690 8700 6780
rect 8550 6600 8730 6690
rect 8580 6510 8760 6600
rect 8610 6480 8760 6510
rect 7530 6360 7680 6420
rect 8610 6390 8790 6480
rect 7500 6300 7680 6360
rect 8640 6300 8820 6390
rect 7500 6270 7650 6300
rect 7470 6210 7650 6270
rect 8670 6270 8820 6300
rect 5940 6120 6090 6210
rect 7440 6150 7620 6210
rect 8670 6150 8850 6270
rect 7410 6120 7620 6150
rect 8700 6120 8850 6150
rect 5940 5940 6120 6120
rect 7410 6090 7590 6120
rect 7380 6060 7560 6090
rect 7350 6030 7560 6060
rect 7320 5970 7530 6030
rect 8700 6000 8880 6120
rect 8730 5970 8880 6000
rect 7290 5940 7500 5970
rect 3600 5910 3870 5940
rect 3540 5880 3900 5910
rect 3510 5850 3900 5880
rect 3450 5820 3900 5850
rect 3420 5790 3900 5820
rect 3360 5760 3900 5790
rect 3300 5730 3900 5760
rect 3270 5700 3900 5730
rect 3210 5670 3900 5700
rect 3180 5640 3900 5670
rect 3120 5610 3900 5640
rect 3090 5580 3530 5610
rect 3030 5550 3480 5580
rect 3000 5520 3450 5550
rect 3000 5490 3390 5520
rect 3000 5460 3330 5490
rect 1590 5430 1830 5460
rect 1560 5310 1830 5430
rect 3000 5430 3300 5460
rect 3000 5400 3240 5430
rect 3000 5370 3180 5400
rect 3000 5340 3150 5370
rect 3000 5310 3090 5340
rect 1560 4710 1860 5310
rect 900 4620 2520 4710
rect 870 4560 2520 4620
rect 900 4470 2520 4560
rect 960 4440 2460 4470
rect 1560 4200 1860 4440
rect 1560 3750 1830 4200
rect 3570 3780 3900 5610
rect 5970 5790 6120 5940
rect 7260 5910 7470 5940
rect 7230 5880 7440 5910
rect 7170 5850 7440 5880
rect 7140 5820 7410 5850
rect 8730 5820 8910 5970
rect 7080 5790 7380 5820
rect 8760 5790 8910 5820
rect 5970 5460 6150 5790
rect 7020 5760 7350 5790
rect 6960 5730 7320 5760
rect 6900 5700 7260 5730
rect 6810 5670 7230 5700
rect 6720 5640 7170 5670
rect 6630 5610 7110 5640
rect 8760 5610 8940 5790
rect 6570 5580 7050 5610
rect 6510 5550 6990 5580
rect 8790 5550 8940 5610
rect 6480 5520 6900 5550
rect 6420 5490 6810 5520
rect 7140 5490 7380 5520
rect 6390 5460 6720 5490
rect 7050 5460 7470 5490
rect 5970 5220 6120 5460
rect 6360 5430 6660 5460
rect 6990 5430 7530 5460
rect 6330 5400 6600 5430
rect 6960 5400 7560 5430
rect 6300 5370 6570 5400
rect 6930 5370 7590 5400
rect 6270 5340 6510 5370
rect 6870 5340 7620 5370
rect 8790 5340 8970 5550
rect 6240 5310 6480 5340
rect 6840 5310 7650 5340
rect 6210 5280 6450 5310
rect 6810 5280 7680 5310
rect 6180 5250 6420 5280
rect 6810 5250 7350 5280
rect 7470 5250 7710 5280
rect 8820 5250 8970 5340
rect 6150 5220 6360 5250
rect 6780 5220 7290 5250
rect 7530 5220 7740 5250
rect 5970 5190 6330 5220
rect 6750 5190 7230 5220
rect 7560 5190 7740 5220
rect 5970 5160 6300 5190
rect 6720 5160 7230 5190
rect 7590 5160 7770 5190
rect 5940 5130 6270 5160
rect 6720 5130 7200 5160
rect 7620 5130 7800 5160
rect 5940 5070 6240 5130
rect 6690 5070 7200 5130
rect 7650 5100 7800 5130
rect 7650 5070 7830 5100
rect 5940 5040 6210 5070
rect 5940 5010 6180 5040
rect 6660 5010 7200 5070
rect 7680 5010 7830 5070
rect 8820 5040 9000 5250
rect 5910 4980 6180 5010
rect 5910 4950 6150 4980
rect 6630 4950 7200 5010
rect 5910 4890 6120 4950
rect 6600 4920 7200 4950
rect 7710 4920 7860 5010
rect 8850 4920 9000 5040
rect 11070 5010 11190 5040
rect 11070 4980 11280 5010
rect 11040 4950 11370 4980
rect 11040 4920 11400 4950
rect 5880 4830 6090 4890
rect 6600 4860 7230 4920
rect 7710 4890 7890 4920
rect 7680 4860 7890 4890
rect 6570 4830 7260 4860
rect 7650 4830 7890 4860
rect 5880 4770 6060 4830
rect 6570 4800 7320 4830
rect 7620 4800 7890 4830
rect 6570 4770 7410 4800
rect 7530 4770 7890 4800
rect 5850 4740 6030 4770
rect 5880 4710 6030 4740
rect 5880 4680 6000 4710
rect 6570 4500 7890 4770
rect 8850 4740 9030 4920
rect 11070 4890 11460 4920
rect 11100 4860 11490 4890
rect 11220 4830 11520 4860
rect 11280 4800 11520 4830
rect 11340 4770 11550 4800
rect 11370 4740 11550 4770
rect 8880 4710 9030 4740
rect 8880 4650 9060 4710
rect 11400 4680 11580 4740
rect 8880 4620 9090 4650
rect 11430 4620 11580 4680
rect 8910 4590 9090 4620
rect 10920 4590 11040 4620
rect 8910 4560 9120 4590
rect 8940 4500 9120 4560
rect 10890 4530 11070 4590
rect 10860 4500 11070 4530
rect 6600 4410 7890 4500
rect 8970 4410 9150 4500
rect 6630 4320 7860 4410
rect 6660 4290 7860 4320
rect 9000 4350 9150 4410
rect 10860 4380 11040 4500
rect 11430 4470 11610 4620
rect 11430 4440 11640 4470
rect 11460 4410 11640 4440
rect 11460 4380 11670 4410
rect 10800 4350 11040 4380
rect 11490 4350 11670 4380
rect 6660 4260 7830 4290
rect 6690 4230 7830 4260
rect 6720 4200 7830 4230
rect 9000 4200 9180 4350
rect 10770 4320 11040 4350
rect 10740 4290 11010 4320
rect 11520 4290 11700 4350
rect 10710 4260 10950 4290
rect 10680 4230 10920 4260
rect 6720 4170 7800 4200
rect 6750 4140 7800 4170
rect 9030 4140 9180 4200
rect 10650 4200 10890 4230
rect 10650 4170 10830 4200
rect 10620 4140 10800 4170
rect 6780 4110 7770 4140
rect 6810 4080 7770 4110
rect 6840 4050 7740 4080
rect 6840 4020 7710 4050
rect 6870 3990 7710 4020
rect 6930 3960 7680 3990
rect 9030 3960 9210 4140
rect 10590 4110 10800 4140
rect 11550 4110 11730 4290
rect 10590 4080 10770 4110
rect 11520 4080 11730 4110
rect 10590 4050 10740 4080
rect 11520 4050 11700 4080
rect 6960 3930 7650 3960
rect 6990 3900 7590 3930
rect 9060 3900 9210 3960
rect 10560 3990 10740 4050
rect 11490 4020 11700 4050
rect 11460 3990 11670 4020
rect 7050 3870 7560 3900
rect 7110 3840 7500 3870
rect 7230 3810 7320 3840
rect 3060 3750 4350 3780
rect 9060 3750 9240 3900
rect 1590 3720 1830 3750
rect 3030 3720 4380 3750
rect 3000 3690 4380 3720
rect 9090 3690 9240 3750
rect 10560 3840 10710 3990
rect 11400 3960 11640 3990
rect 11370 3930 11640 3960
rect 11310 3900 11580 3930
rect 11250 3870 11550 3900
rect 11220 3840 11520 3870
rect 10560 3720 10740 3840
rect 11220 3810 11460 3840
rect 11220 3780 11430 3810
rect 11250 3750 11460 3780
rect 10590 3690 10770 3720
rect 11280 3690 11490 3750
rect 3000 3600 4410 3690
rect 3000 3540 4380 3600
rect 9090 3570 9270 3690
rect 10590 3660 10800 3690
rect 11310 3660 11520 3690
rect 10620 3630 10830 3660
rect 11340 3630 11550 3660
rect 10620 3600 10860 3630
rect 11370 3600 11550 3630
rect 10650 3570 10860 3600
rect 3030 3510 4380 3540
rect 9120 3540 9270 3570
rect 10620 3540 10860 3570
rect 11400 3540 11580 3600
rect 9120 3450 9300 3540
rect 10590 3510 10860 3540
rect 10560 3480 10800 3510
rect 10560 3450 10770 3480
rect 5940 3390 6000 3420
rect 5910 3360 6030 3390
rect 9150 3360 9330 3450
rect 10530 3420 10740 3450
rect 10530 3390 10710 3420
rect 10500 3360 10710 3390
rect 5880 3330 6060 3360
rect 5850 3270 6060 3330
rect 9180 3270 9360 3360
rect 10500 3300 10680 3360
rect 11430 3330 11610 3540
rect 11400 3300 11580 3330
rect 5820 3240 6030 3270
rect 5790 3210 6000 3240
rect 9210 3210 9390 3270
rect 5790 3180 5970 3210
rect 5760 3150 5970 3180
rect 9240 3150 9420 3210
rect 5760 3120 5940 3150
rect 9240 3120 9450 3150
rect 5730 3090 5940 3120
rect 9270 3090 9450 3120
rect 10500 3120 10650 3300
rect 11370 3240 11580 3300
rect 11340 3210 11550 3240
rect 11310 3180 11520 3210
rect 11250 3150 11520 3180
rect 11220 3120 11490 3150
rect 5730 3060 5910 3090
rect 9270 3060 9480 3090
rect 5700 2970 5880 3060
rect 9300 3030 9480 3060
rect 9300 3000 9510 3030
rect 10500 3000 10680 3120
rect 11220 3090 11460 3120
rect 11190 3060 11430 3090
rect 11220 3030 11370 3060
rect 11250 3000 11340 3030
rect 9330 2970 9540 3000
rect 10530 2970 10710 3000
rect 5670 2880 5850 2970
rect 9360 2940 9570 2970
rect 10530 2940 10740 2970
rect 9360 2910 9600 2940
rect 10560 2910 10770 2940
rect 9390 2880 9660 2910
rect 10560 2880 10800 2910
rect 5670 2850 5820 2880
rect 5640 2670 5820 2850
rect 9420 2850 9720 2880
rect 10590 2850 10830 2880
rect 9420 2820 9840 2850
rect 10620 2820 10890 2850
rect 9450 2790 9960 2820
rect 10650 2790 10950 2820
rect 9510 2760 10050 2790
rect 10680 2760 10980 2790
rect 9570 2730 10170 2760
rect 10710 2730 10980 2760
rect 9630 2700 10230 2730
rect 10740 2700 10980 2730
rect 9720 2670 10290 2700
rect 10800 2670 10950 2700
rect 5670 2640 5820 2670
rect 9870 2640 10350 2670
rect 10860 2640 10920 2670
rect 5670 2550 5850 2640
rect 9960 2610 10410 2640
rect 10050 2580 10440 2610
rect 10140 2550 10470 2580
rect 5700 2520 5880 2550
rect 10230 2520 10530 2550
rect 5700 2490 5910 2520
rect 10290 2490 10560 2520
rect 5730 2460 5910 2490
rect 10320 2460 10590 2490
rect 5730 2430 5940 2460
rect 10380 2430 10620 2460
rect 5700 2400 5970 2430
rect 10410 2400 10650 2430
rect 5670 2370 6000 2400
rect 10440 2370 10680 2400
rect 5610 2340 6030 2370
rect 10470 2340 10710 2370
rect 5580 2310 6060 2340
rect 10500 2310 10710 2340
rect 5520 2280 5820 2310
rect 5850 2280 6120 2310
rect 10530 2280 10740 2310
rect 5490 2250 5790 2280
rect 5880 2250 6180 2280
rect 7290 2250 7350 2280
rect 5430 2220 5760 2250
rect 5910 2220 6240 2250
rect 7260 2220 7380 2250
rect 10560 2220 10770 2280
rect 5400 2190 5700 2220
rect 5970 2190 6300 2220
rect 7230 2190 7410 2220
rect 10590 2190 10800 2220
rect 5370 2160 5640 2190
rect 6000 2160 6390 2190
rect 7200 2160 7410 2190
rect 5340 2130 5610 2160
rect 6030 2130 6450 2160
rect 7140 2130 7410 2160
rect 10200 2130 10260 2160
rect 10620 2130 10800 2190
rect 5280 2100 5580 2130
rect 6090 2100 6570 2130
rect 7080 2100 7380 2130
rect 5280 2070 5520 2100
rect 6150 2070 6810 2100
rect 6960 2070 7350 2100
rect 10170 2070 10320 2130
rect 5250 2040 5490 2070
rect 6210 2040 7320 2070
rect 5250 2010 5460 2040
rect 6270 2010 7260 2040
rect 5250 1980 5400 2010
rect 6360 1980 7200 2010
rect 5250 1950 5370 1980
rect 6450 1950 7140 1980
rect 5250 1920 5340 1950
rect 6600 1920 7050 1950
rect 5250 1890 5310 1920
rect 6810 1890 7050 1920
rect 10140 1920 10320 2070
rect 10650 2040 10830 2130
rect 10680 2010 10830 2040
rect 10140 1890 10290 1920
rect 5250 1860 5280 1890
rect 6840 1860 7080 1890
rect 10110 1860 10290 1890
rect 6870 1830 7110 1860
rect 10080 1830 10290 1860
rect 6870 1800 7140 1830
rect 6900 1770 7170 1800
rect 10050 1770 10260 1830
rect 10680 1800 10860 2010
rect 6930 1740 7200 1770
rect 10050 1740 10230 1770
rect 10680 1740 10830 1800
rect 6960 1710 7230 1740
rect 8820 1710 8880 1740
rect 10080 1710 10200 1740
rect 6990 1680 7260 1710
rect 8790 1680 8940 1710
rect 10110 1680 10170 1710
rect 7020 1650 7290 1680
rect 8790 1650 8970 1680
rect 7050 1620 7350 1650
rect 8760 1620 9000 1650
rect 10650 1620 10830 1740
rect 7080 1590 7380 1620
rect 8790 1590 9060 1620
rect 7140 1560 7410 1590
rect 8820 1560 9090 1590
rect 7170 1530 7470 1560
rect 8850 1530 9120 1560
rect 10620 1530 10800 1620
rect 7200 1500 7530 1530
rect 8880 1500 9150 1530
rect 7260 1470 7560 1500
rect 8910 1470 9180 1500
rect 10590 1470 10770 1530
rect 7290 1440 7620 1470
rect 8970 1440 9240 1470
rect 10560 1440 10770 1470
rect 7350 1410 7680 1440
rect 9000 1410 9270 1440
rect 10560 1410 10740 1440
rect 7380 1380 7710 1410
rect 9030 1380 9300 1410
rect 10530 1380 10740 1410
rect 7440 1350 7770 1380
rect 9090 1350 9330 1380
rect 10530 1350 10710 1380
rect 7470 1320 7830 1350
rect 9120 1320 9360 1350
rect 10500 1320 10710 1350
rect 7530 1290 7890 1320
rect 9150 1290 9420 1320
rect 10470 1290 10680 1320
rect 7590 1260 7950 1290
rect 9180 1260 9450 1290
rect 10470 1260 10650 1290
rect 7650 1230 7980 1260
rect 9210 1230 9480 1260
rect 10440 1230 10650 1260
rect 7680 1200 8040 1230
rect 9270 1200 9510 1230
rect 10410 1200 10620 1230
rect 7740 1170 8100 1200
rect 9300 1170 9540 1200
rect 10380 1170 10590 1200
rect 7800 1140 8190 1170
rect 9330 1140 9600 1170
rect 10350 1140 10590 1170
rect 7860 1110 8250 1140
rect 9360 1110 9630 1140
rect 10350 1110 10560 1140
rect 7920 1080 8340 1110
rect 9390 1080 9660 1110
rect 10320 1080 10530 1110
rect 7980 1050 8400 1080
rect 9420 1050 9690 1080
rect 10290 1050 10500 1080
rect 8040 1020 8490 1050
rect 9420 1020 9750 1050
rect 10260 1020 10470 1050
rect 8100 990 8580 1020
rect 9360 990 9780 1020
rect 10230 990 10440 1020
rect 8160 960 8700 990
rect 9300 960 9840 990
rect 10200 960 10440 990
rect 8220 930 8910 960
rect 9150 930 9540 960
rect 9600 930 9900 960
rect 10170 930 10410 960
rect 8310 900 9510 930
rect 9630 900 9960 930
rect 10110 900 10380 930
rect 8370 870 9480 900
rect 9690 870 10020 900
rect 10080 870 10350 900
rect 8460 840 9420 870
rect 9720 840 10320 870
rect 8580 810 9360 840
rect 9780 810 10260 840
rect 8700 780 9300 810
rect 9810 780 10230 810
rect 8970 750 9060 780
rect 9870 750 10200 780
rect 9930 720 10170 750
<< end >>
